typedef uvm_sequencer#(read_tx) read_sqr;
